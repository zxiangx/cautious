/******************************************************************************
 ** Logisim goes FPGA automatic generated Verilog code                       **
 **                                                                          **
 ** Component : RegFile                                                      **
 **                                                                          **
 ******************************************************************************/

`timescale 1ns/1ps
module RegFile( Clk,
                Din,
                R1Adr,
                R2Adr,
                WAdr,
                WE,
                R1,
                R2);

   /***************************************************************************
    ** Here the inputs are defined                                           **
    ***************************************************************************/
   input  Clk;
   input[31:0]  Din;
   input[4:0]  WAdr;
   input  WE;
   input[4:0]  R1Adr;
   input[4:0]  R2Adr;

   /***************************************************************************
    ** Here the outputs are defined                                          **
    ***************************************************************************/
   output reg[31:0] R1;
   output reg[31:0] R2;

   /***************************************************************************
    ** Internal register file definition                                     **
    ***************************************************************************/
   reg[31:0] reg_file[31:0]; // 32�?32位的寄存�?

   integer i;

   // 初始化寄存器文件（可选）
   initial begin
      for (i = 0; i < 32; i = i + 1) begin
         reg_file[i] = 32'b0;
      end
   end

   /***************************************************************************
    ** Write operation                                                       **
    ***************************************************************************/
   always @(posedge Clk) begin
      if (WE) begin
         // 写操作，WE为高电平时写入数�?
         reg_file[WAdr] <= Din;
      end
   end

   /***************************************************************************
    ** Read operation                                                        **
    ***************************************************************************/
   always @(*) begin
      // 读操作：根据输入的寄存器编号读取寄存器文件中的数�?
      R1 = reg_file[R1Adr];
      R2 = reg_file[R2Adr];
   end

endmodule
